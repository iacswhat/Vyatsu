// megafunction wizard: %LPM_CLSHIFT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_clshift 

// ============================================================
// File Name: RG3S.v
// Megafunction Name(s):
// 			lpm_clshift
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module RG3S (
	data,
	direction,
	distance,
	result);

	input	[46:0]  data;
	input	  direction;
	input	  distance;
	output	[46:0]  result;

	wire [46:0] sub_wire0;
	wire [46:0] result = sub_wire0[46:0];
	wire  sub_wire1 = distance;
	wire  sub_wire2 = sub_wire1;

	lpm_clshift	lpm_clshift_component (
				.distance (sub_wire2),
				.direction (direction),
				.data (data),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock (),
				.overflow (),
				.underflow ()
				// synopsys translate_on
				);
	defparam
		lpm_clshift_component.lpm_shifttype = "LOGICAL",
		lpm_clshift_component.lpm_type = "LPM_CLSHIFT",
		lpm_clshift_component.lpm_width = 47,
		lpm_clshift_component.lpm_widthdist = 1;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: LPM_SHIFTTYPE NUMERIC "0"
// Retrieval info: PRIVATE: LPM_WIDTH NUMERIC "47"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: lpm_width_varies NUMERIC "0"
// Retrieval info: PRIVATE: lpm_widthdist NUMERIC "1"
// Retrieval info: PRIVATE: lpm_widthdist_style NUMERIC "1"
// Retrieval info: PRIVATE: port_direction NUMERIC "2"
// Retrieval info: CONSTANT: LPM_SHIFTTYPE STRING "LOGICAL"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_CLSHIFT"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "47"
// Retrieval info: CONSTANT: LPM_WIDTHDIST NUMERIC "1"
// Retrieval info: USED_PORT: data 0 0 47 0 INPUT NODEFVAL data[46..0]
// Retrieval info: USED_PORT: direction 0 0 0 0 INPUT NODEFVAL direction
// Retrieval info: USED_PORT: distance 0 0 0 0 INPUT NODEFVAL distance
// Retrieval info: USED_PORT: result 0 0 47 0 OUTPUT NODEFVAL result[46..0]
// Retrieval info: CONNECT: @distance 0 0 1 0 distance 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 47 0 data 0 0 47 0
// Retrieval info: CONNECT: result 0 0 47 0 @result 0 0 47 0
// Retrieval info: CONNECT: @direction 0 0 0 0 direction 0 0 0 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL RG3S.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL RG3S.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL RG3S.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL RG3S.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL RG3S_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL RG3S_bb.v TRUE
